library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity rom is
   port( clk      : in std_logic;
         endereco : in unsigned(6 downto 0);
         dado     : out unsigned(16 downto 0) 
   );
end entity;
architecture a_rom of rom is
   type mem is array (0 to 127) of unsigned(16 downto 0);
   constant conteudo_rom : mem := (
      -- caso endereco => conteudo
      0  => B"0011_0001110_1000_10", -- ld 14 into accumulator
      1  => B"0101_0000000_0101_00", -- Accumulator -> r5
      2  => B"0111_0000011_0101_00", -- subi r5, 3
      3  => B"1001_0001011_0101_11", -- cmpi r5, 11
      4  => B"1001_0001010_0000_00", -- cmpi r5, 10
      5  => B"00000000000000101",
      6  => B"0011_0000001_0001_10", -- ld into r1
      7  => B"0011_0100001_0011_10", -- ld into r3
      8  => B"0010_0000000_0011_00", -- add r3
      9  => B"0100_0000000_0001_00", -- sub r1
      10 => B"0101_0000000_1110_10", -- load r6 into Accumulator
      11 => B"11110000000001011", -- B. instruction says "jump to 0"
      -- abaixo: casos omissos => (zero em todos os bits)
      others => (others=>'0')
   );
begin
   process(clk)
   begin
      if(rising_edge(clk)) then
         dado <= conteudo_rom(to_integer(endereco));
      end if;
   end process;
end architecture;