library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity rom is
   port( clk      : in std_logic;
         endereco : in unsigned(6 downto 0);
         dado     : out unsigned(16 downto 0) 
   );
end entity;
architecture a_rom of rom is
   type mem is array (0 to 127) of unsigned(16 downto 0);
   constant conteudo_rom : mem := ( 
      -- load data into RAM     
      0  => B"0011_0000000_1000_00", -- ld A,0
      -- R3 += 1
      1  => B"0101_0000000_1011_00", -- mv A,R3
      2  => B"0110_0000001_0100_00", -- addi 1
      3  => B"0101_0000000_0011_00", -- mv R3,A
      -- SW R3 into address R3
      4  => B"1110_0000001_0011_00", -- SW R3
      -- Repeat 32 times
      5  => B"0111_0100000_0000_00", -- subi 32  
      6  => B"1101_1111011_0000_00", -- BMI -5 0000101 1111011 

      -- Remove multiples of 2
      7  => B"0011_0000000_1000_00", -- ld A,0
      -- R4 += 2
      8  => B"0101_0000000_1100_00", -- mv A,R4
      9  => B"0110_0000010_0100_00", -- addi 2
      10 => B"0101_0000000_0100_00", -- mv R4,A
      -- SW 0 into address R4
      11 => B"1000_0000000_1000_00", -- clr A
      12 => B"1110_0000001_0100_00", -- SW R4
      13 => B"0101_0000000_1100_00", -- mv A,R4
      14 => B"0111_0100000_0000_00", -- subi 32  
      15 => B"1101_1111001_0000_00", -- BMI -7 0000111 1111000 1111001

      -- Remove multiples of 3
      -- reset accumulator and R4
      16 => B"0011_0000000_1000_00", -- ld A,0
      17 => B"0101_0000000_0100_00", -- mv R4,A
      -- R4 += 3
      18 => B"0101_0000000_1100_00", -- mv A,R4
      19 => B"0110_0000011_0100_00", -- addi 3
      20 => B"0101_0000000_0100_00", -- mv R4,A
      -- SW 0 into address R4
      21 => B"1000_0000000_1000_00", -- clr A
      22 => B"1110_0000001_0100_00", -- SW R4
      23 => B"0101_0000000_1100_00", -- mv A,R4
      24 => B"0111_0100000_0000_00", -- subi 32  
      25 => B"1101_1111001_0000_00", -- BMI -7 0000111 1111000 1111001

      -- Remove multiples of 5
      -- reset accumulator and R4
      26 => B"0011_0000000_1000_00", -- ld A,0
      27 => B"0101_0000000_0100_00", -- mv R4,A
      -- R4 += 5
      28 => B"0101_0000000_1100_00", -- mv A,R4
      29 => B"0110_0000101_0100_00", -- addi 5
      30 => B"0101_0000000_0100_00", -- mv R4,A
      -- SW 0 into address R4
      31 => B"1000_0000000_1000_00", -- clr A
      32 => B"1110_0000001_0100_00", -- SW R4
      33 => B"0101_0000000_1100_00", -- mv A,R4
      34 => B"0111_0100000_0000_00", -- subi 32  
      35 => B"1101_1111001_0000_00", -- BMI -7 0000111 1111000 1111001

      -- write prime numbers into R0
      -- accumulator and R3 <= 1
      36 => B"0011_0000001_1000_00", -- ld A,1
      37 => B"0101_0000000_0011_00", -- mv R3,A
      -- R3 += 1
      38 => B"0101_0000000_1011_00", -- mv A,R3
      39 => B"0110_0000001_0100_00", -- addi 1
      40 => B"0101_0000000_0011_00", -- mv R3,A
      -- LW R3
      41 => B"1110_0000001_0011_01", -- LW R3
      -- Write R3 into R0
      42 => B"0101_0000000_0000_00", -- mv R0,A
      -- Repeat 32 times
      43 => B"0111_0011111_0000_00", -- subi 31  0011111
      44 => B"1101_1111010_0000_00", -- BMI -6 0000110 1111001 1111010




      --0  => B"0011_0001010_1000_00", -- ld A,10
     --1  => B"0101_0000000_0011_00", -- mv R3,A
     -- 2  => B"0101_0000000_0100_00", -- mv R4,A
     -- 3  => B"0011_0011001_1000_00", -- ld A,25
      --4  => B"1110_0000001_0011_00", -- SW R3
      --5  => B"1000_0000000_1000_00", -- clr A
      --6  => B"1110_0000001_0011_01", -- LW R3
      



      --1  => B"0011_0000101_0100_00", -- ld R4,5
      --2  => B"0010_0000000_0011_00", -- add A,R3
      --4  => B"0100_0000000_0100_00", -- sub A,R4
      --5  => B"0110_0010001_0100_00", -- addi 17
      --6  => B"0110_1111011_0011_00", -- addi -5 
      --7  => B"0111_0001010_0000_00", -- subi 10
      --8  => B"1010_1111000_0000_00", -- BEQ -8

      --0  => B"0011_0000101_0011_10", -- ld R3,5
      --1  => B"0011_0001000_0100_00", -- ld R4,8
      --2  => B"0010_0000000_0011_00", -- add A,R3
      --3  => B"0010_0000000_0100_00", -- add A,R4
      --4  => B"0101_0000000_0101_00", -- mv R5,A
      --5  => B"0111_0000001_0101_00", -- subi 1,R5
      --6  => B"1111_0010100_0000_00", -- j 20
      --7  => B"1000_0000000_0101_00", -- clr R5

      --20 => B"0101_0000000_1101_00", -- mv A,R5
      --21 => B"0101_0000000_0011_00", -- mv R3,A
      --22 => B"1111_0000010_0000_00", -- j 2
      --23  => B"1000_0000000_0011_00", -- clr R3

      -- caso endereco => conteudo
      --0  => B"0011_0001110_1000_10", -- ld 14 into accumulator
      --1  => B"0101_0000000_0101_00", -- MOV Accumulator -> r5
      --2  => B"0111_0000011_0101_00", -- subi r5, 3
      --3  => B"1001_0001011_0101_11", -- cmpi r5, 11
      --4  => B"1001_0001010_0000_00", -- cmpi r5, 10
      --5  => B"0111_0001001_0101_01", -- subi r5, 9
      --6  => B"0011_0000001_0001_10", -- ld into r1
      --7  => B"0011_0100001_0011_10", -- ld into r3
      --8  => B"0010_0000000_0011_00", -- add r3
      --9  => B"0100_0000000_0001_00", -- sub r1
      --10 => B"0101_0000000_1110_10", -- load r6 into Accumulator
      --11 => B"11110000000001011", -- B. instruction says "jump to 0"
      -- abaixo: casos omissos => (zero em todos os bits)
      others => (others=>'0')
   );
begin
   process(clk)
   begin
      if(rising_edge(clk)) then
         dado <= conteudo_rom(to_integer(endereco));
      end if;
   end process;
end architecture;