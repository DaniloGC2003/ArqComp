library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity rom is
   port( clk      : in std_logic;
         endereco : in unsigned(6 downto 0);
         dado     : out unsigned(16 downto 0) 
   );
end entity;
architecture a_rom of rom is
   type mem is array (0 to 127) of unsigned(16 downto 0);
   constant conteudo_rom : mem := ( 
      -- R2: stores the current value to be used in the RAM
      -- R3: stores the current address to be used in the RAM

      -- R0: iterator
         0  => B"0011_0100000_1000_00", -- ld A,32
         1  => B"0101_0000000_0000_00", -- mv R0,A
      -- R1: address and data to be used in RAM
         2  => B"0011_0000001_1000_00", -- ld A,1
         3  => B"0101_0000000_0001_00", -- mv R1,A

      -- Fill up RAM addrs 1 to 32
         -- Store R1 in R1
            4  => B"1110_0000001_0001_00", -- SW R1,R1
         -- R1 += 1
            5  => B"0101_0000000_1001_00", -- mv A,R1
            6  => B"0110_0000001_0100_00", -- addi 1
            7  => B"0101_0000000_0001_00", -- mv R1,A
         -- DJNZ 4,R4
            8  => B"0001_0000100_0000_00", -- DJNZ 4,R0

      -- Remove multiples of 2
         -- clear A and R4
            9  => B"1000_0000000_1000_00", -- clr A
            10 => B"0101_0000000_0100_00", -- mv R4,A
         -- R0 <= 16 (loop will be executed 16 times)
            11  => B"0011_0010000_1000_00", -- ld A,16
            12  => B"0101_0000000_0000_00", -- mv R0,A 
         -- R4 += 2
            13  => B"0101_0000000_1100_00", -- mv A,R4
            14  => B"0110_0000010_0100_00", -- addi 2
            15 => B"0101_0000000_0100_00", -- mv R4,A
         -- SW R2 (storing 0) into address R4
            16  => B"1110_0000010_0100_00", -- SW R2,R4
            --17 => B"0101_0000000_1100_00", -- mv A,R4
         -- DJNZ 13,R0
            17  => B"0001_0001101_0000_00", -- DJNZ 13,R0





                     -- R0 -= 1 (so that, at the end of the loop, R0 is decremented by 2)
            --16  => B"0101_0000000_1000_00", -- mv A,R0
            --17  => B"0111_0000001_0000_00", -- subi 1
            --18 => B"0101_0000000_0000_00", -- mv R0,A


      -- Remove multiples of 2
         -- Reset iterator R4
            -- A = 64
               --26  => B"0011_0100000_1000_00", -- ld A,32
               --27  => B"0110_0100000_0100_00", -- addi 32
               --28  => B"0110_0100000_0100_00", -- addi 32
               --29  => B"0110_0100000_0100_00", -- addi 32
            -- R4 = 128
               --30  => B"0101_0000000_0100_00", -- mv R4,A
         -- clear A, R2 and R3
            --31  => B"1000_0000000_1000_00", -- clr A
            --32  => B"0101_0000000_0010_00", -- mv R2,A
            --33  => B"0101_0000000_0011_00", -- mv R3,A
         -- R5 reads data in address R3
            --34  => B"1110_0000101_0011_01", -- LW R5,R3
         -- keep subtracting 2 from R5 until it's equal to 0 (in this case, it's a multiple of 2) or negative 
         -- RESULTADO NEGATIVO: AINDA N SEI; RESULTADO 0: MULTIPLO DE 2; RESULTADO POSITIVO: NAO É MULTIPLO DE 2
         -- Clear R1
            --35  => B"1000_0000000_1000_00", -- clr A
            --36  => B"0101_0000000_0001_00", -- mv R1,A
         -- R1 += 2
            --35  => B"0101_0000000_1001_00", -- mv A,R1
            --36  => B"0110_0000010_0100_00", -- addi 2       A = 2          A
            --37  => B"0101_0000000_0001_00", -- mv R1,A  
         -- check if result is positive, negative or zero
            --38  => B"0100_0000000_0101_00", -- sub A,R5    
            --39  => B"1101_1111100_0000_00", -- BMI -4
         -- check if result is zero. If so, remove from RAM
         --30  => B"0101_0000000_1101_00", -- mv A,R5
         --79  => B"0111_0000010_0000_00", -- subi 2

         -- Store 0 in R3
         --29  => B"1110_0000010_0011_00", -- SW R2,R3
         -- R3 += 1
            --40  => B"0101_0000000_1011_00", -- mv A,R3
            --41  => B"0110_0000001_0100_00", -- addi 1
            --42  => B"0101_0000000_0011_00", -- mv R3,A
         -- DJNZ 15,R4
            --43  => B"0001_0100010_0100_00", -- DJNZ 34,R4 0100010


      --1  => B"0101_0000000_0001_00", -- mv R1,A
      --3  => B"0001_0000010_0001_00", -- DJNZ 2,R1

      --0  => B"0011_0100001_1000_00", -- ld A,33
      --1  => B"0101_0000000_0001_00", -- mv R1,A
      --2  => B"0011_0000101_1000_00", -- ld A,5
      --3  => B"0101_0000000_0000_00", -- mv R0,A
      --4  => B"0100_0000000_0000_00", -- sub A,R0
      --5  => B"0001_0001110_0001_00", -- DJNZ 14,R1
      --6  => B"0011_0001010_1000_00", -- ld A,10
      --7  => B"0100_0000000_0000_00", -- sub A,R0
      --8  => B"0001_0001110_0001_00", -- DJNZ 14,R1

   

      


      --0  => B"0011_0001010_1000_00", -- ld A,10
     --1  => B"0101_0000000_0011_00", -- mv R3,A
     -- 2  => B"0101_0000000_0100_00", -- mv R4,A
     -- 3  => B"0011_0011001_1000_00", -- ld A,25
      --4  => B"1110_0000001_0011_00", -- SW R3
      --5  => B"1000_0000000_1000_00", -- clr A
      --6  => B"1110_0000001_0011_01", -- LW R3
      



      --1  => B"0011_0000101_0100_00", -- ld R4,5
      --2  => B"0010_0000000_0011_00", -- add A,R3
      --4  => B"0100_0000000_0100_00", -- sub A,R4
      --5  => B"0110_0010001_0100_00", -- addi 17
      --6  => B"0110_1111011_0011_00", -- addi -5 
      --7  => B"0111_0001010_0000_00", -- subi 10
      --8  => B"1010_1111000_0000_00", -- BEQ -8

      --0  => B"0011_0000101_0011_10", -- ld R3,5
      --1  => B"0011_0001000_0100_00", -- ld R4,8
      --2  => B"0010_0000000_0011_00", -- add A,R3
      --3  => B"0010_0000000_0100_00", -- add A,R4
      --4  => B"0101_0000000_0101_00", -- mv R5,A
      --5  => B"0111_0000001_0101_00", -- subi 1,R5
      --6  => B"1111_0010100_0000_00", -- j 20
      --7  => B"1000_0000000_0101_00", -- clr R5

      --20 => B"0101_0000000_1101_00", -- mv A,R5
      --21 => B"0101_0000000_0011_00", -- mv R3,A
      --22 => B"1111_0000010_0000_00", -- j 2
      --23  => B"1000_0000000_0011_00", -- clr R3

      -- caso endereco => conteudo
      --0  => B"0011_0001110_1000_10", -- ld 14 into accumulator
      --1  => B"0101_0000000_0101_00", -- MOV Accumulator -> r5
      --2  => B"0111_0000011_0101_00", -- subi r5, 3
      --3  => B"1001_0001011_0101_11", -- cmpi r5, 11
      --4  => B"1001_0001010_0000_00", -- cmpi r5, 10
      --5  => B"0111_0001001_0101_01", -- subi r5, 9
      --6  => B"0011_0000001_0001_10", -- ld into r1
      --7  => B"0011_0100001_0011_10", -- ld into r3
      --8  => B"0010_0000000_0011_00", -- add r3
      --9  => B"0100_0000000_0001_00", -- sub r1
      --10 => B"0101_0000000_1110_10", -- load r6 into Accumulator
      --11 => B"11110000000001011", -- B. instruction says "jump to 0"
      -- abaixo: casos omissos => (zero em todos os bits)
      others => (others=>'0')
   );
begin
   process(clk)
   begin
      if(rising_edge(clk)) then
         dado <= conteudo_rom(to_integer(endereco));
      end if;
   end process;
end architecture;